module mant_normaliser
(
    input wire [48:0] pre_res_mant,
    input wire [7:0] exp_max,
    
    output wire []
)

endmodule